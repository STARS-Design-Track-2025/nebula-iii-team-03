`default_nettype none
module player_lut #(parameter int player_height = 20, parameter int player_width = 15)
(   
    //[0:11] Means you have 12 characters. Alaphabet input is 5 bits and gives you acces to 2^6 characters!!
    input logic [3:0] player_state,
    input logic is_1_displayed, p1Left, p2Left,
    input logic is_2_displayed,
    output logic [(player_height * player_width * 8)-1:0] player
);
     
    logic [299:0][7:0] player_sprite;
    logic [1:0] player_select;
    


    always_comb begin
        player_select = 0;
        if(is_1_displayed) begin
            player_select = player_state[1:0];
        end
        else if(is_2_displayed) begin
            player_select = player_state[3:2];
        end
        else if(is_1_displayed && is_2_displayed) begin
            player_select = player_state[1:0];
        end
        else begin
            player_select  = 0;
        end

        case(player_select) 

        2'd0: begin
         player_sprite[299:285] = {8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000};
         player_sprite[284:270] = {8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000};
         player_sprite[269:255] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000};
         player_sprite[254:240] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000};
         player_sprite[239:225] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[224:210] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[209:195] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[194:180] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11100000};
         player_sprite[179:165] = {8'b00000000, 8'b11111001, 8'b11100000, 8'b01000100, 8'b11100000, 8'b11100000, 8'b11111001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111001, 8'b00000000, 8'b01000100, 8'b11100000, 8'b11100000};
         player_sprite[164:150] = {8'b00000000, 8'b11111001, 8'b11100000, 8'b01000100, 8'b11100000, 8'b11100000, 8'b11111001, 8'b11111001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111001, 8'b01000100, 8'b11100000, 8'b00000000};
         player_sprite[149:135] = {8'b00000000, 8'b11111001, 8'b11111001, 8'b01000100, 8'b11100000, 8'b11100000, 8'b11111001, 8'b11111001, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000};
         player_sprite[134:120] = {8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111111, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000};
         player_sprite[119:105] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11111001, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[104:90] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[89:75] = {8'b00000000, 8'b11100000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[74:60] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b11111001, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[59:45] = {8'b00000000, 8'b00000000, 8'b11100000, 8'b01000100, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[44:30] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[29:15] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[14:0] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        end


        2'd1: begin
         player_sprite[299:285] = {8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[284:270] = {8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[269:255] = {8'b00000000, 8'b11111001, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[254:240] = {8'b00000000, 8'b11111111, 8'b11111111, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[239:225] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[224:210] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[209:195] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[194:180] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b11100000, 8'b11100000, 8'b00000000, 8'b11111111, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[179:165] = {8'b00000000, 8'b00000000, 8'b11111001, 8'b11100000, 8'b11100000, 8'b11111001, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[164:150] = {8'b00000000, 8'b00000000, 8'b11111001, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[149:135] = {8'b00000000, 8'b00000000, 8'b11111001, 8'b01000100, 8'b11111001, 8'b01000100, 8'b01000100, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11111001, 8'b11100000};
         player_sprite[134:120] = {8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11100000, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b11100000};
         player_sprite[119:105] = {8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111111, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11100000, 8'b11100000};
         player_sprite[104:90] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[89:75] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[74:60] = {8'b00000000, 8'b00000000, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b00000000, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[59:45] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b11100000, 8'b00000000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[44:30] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[29:15] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[14:0] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

         end

        2'd2: begin
         player_sprite[299:285] = {8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000};
         player_sprite[284:270] = {8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000};
         player_sprite[269:255] = {8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[254:240] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[239:225] = {8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b01000100, 8'b00000000};
         player_sprite[224:210] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[209:195] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[194:180] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[179:165] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11100000, 8'b11100000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b00000000};
         player_sprite[164:150] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b11100000, 8'b11100000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b00000000};
         player_sprite[149:135] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11111111, 8'b00000000, 8'b11100000, 8'b11100000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b00000000};
         player_sprite[134:120] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[119:105] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111111, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b11100000, 8'b11100000, 8'b00000000};
         player_sprite[104:90] = {8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b00000000, 8'b01000100, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b11100000, 8'b11100000, 8'b00000000};
         player_sprite[89:75] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b11100000, 8'b00000000, 8'b11111001, 8'b00000000, 8'b11111001, 8'b11111001, 8'b11111001, 8'b11111001, 8'b00000000, 8'b00000000, 8'b11100000, 8'b00000000};
         player_sprite[74:60] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[59:45] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b11100000, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[44:30] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000};
         player_sprite[29:15] = {8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b00000000, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000};
         player_sprite[14:0] = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

        
        end
        default: player_sprite = 0;
        endcase
    // player_height = 30, parameter int player_width = 19
    if(is_1_displayed) begin
    if(~p1Left) begin //Regular
    for(int i = 0; i < player_height ; i++) begin
        for(int j = 0; j < player_width; j++) begin
         player[((player_height * player_width * 8)-1) - (i * player_width + j)*8-:8] = player_sprite[i * player_width + (player_width - 1 - j)];
        
            end
        end
    end
    else begin // Reversed
        for(int i = player_height * player_width - 1; i >= 0 ; i--) begin
        player[((player_height * player_width * 8)-1) - i*8-:8] = player_sprite[i];
    end
    end
    end
    else if(is_2_displayed)begin 
        if(~p2Left) begin //Regular
        for(int i = player_height * player_width - 1; i >= 0 ; i--) begin
        player[((player_height * player_width * 8)-1) - i*8-:8] = player_sprite[i];
        end
    end
        else begin
        for(int i = 0; i < player_height ; i++) begin
            for(int j = 0; j < player_width; j++) begin
                player[((player_height * player_width * 8)-1) - (i * player_width + j)*8-:8] = player_sprite[i * player_width + (player_width - 1 - j)];
            end
        end
        end
    end
    else begin
        player = 0;
    end

    end
endmodule


    