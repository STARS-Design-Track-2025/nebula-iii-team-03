`default_nettype none
module t03_player_lut (
	player_state,
	is_1_displayed,
	p1Left,
	p2Left,
	is_2_displayed,
	player
);
	reg _sv2v_0;
	parameter signed [31:0] player_height = 20;
	parameter signed [31:0] player_width = 15;
	input wire [3:0] player_state;
	input wire is_1_displayed;
	input wire p1Left;
	input wire p2Left;
	input wire is_2_displayed;
	output reg [((player_height * player_width) * 8) - 1:0] player;
	reg [2399:0] player_sprite;
	reg [1:0] player_select;
	always @(*) begin
		if (_sv2v_0)
			;
		player_select = 0;
		if (is_1_displayed)
			player_select = player_state[1:0];
		else if (is_2_displayed)
			player_select = player_state[3:2];
		else if (is_1_displayed && is_2_displayed)
			player_select = player_state[1:0];
		else
			player_select = 0;
		case (player_select)
			2'd0: begin
				player_sprite[2280+:120] = 120'b111110011111100111111001111110010000000000000000000000000000000000000000000000001111100111111001111110011111100100000000;
				player_sprite[2160+:120] = 120'b000000001111100111111001111110010000000000000000000000000000000000000000000000001111100111111001111110011111100100000000;
				player_sprite[2040+:120] = 120'b000000000000000011111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000;
				player_sprite[1920+:120] = 120'b000000000000000011111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000;
				player_sprite[1800+:120] = 120'b000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000;
				player_sprite[1680+:120] = 120'b000000000000000011111111111111111111111100000000111111111111111111111111111111111111111100000000000000000000000000000000;
				player_sprite[1560+:120] = 120'b000000000000000000000000111111111111111111111111000000000000000011111111111111111111111100000000000000000000000000000000;
				player_sprite[1440+:120] = 120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110011111100111100000;
				player_sprite[1320+:120] = 120'b000000001111100111100000010001001110000011100000111110011111111111111111111111111111100100000000010001001110000011100000;
				player_sprite[1200+:120] = 120'b000000001111100111100000010001001110000011100000111110011111100111111111111111111111111111111001010001001110000000000000;
				player_sprite[1080+:120] = 120'b000000001111100111111001010001001110000011100000111110011111100111111111111111111111111111111001111110010000000000000000;
				player_sprite[960+:120] = 120'b000000000000000011111001111110011111111111111001111110010000000000000000111111111111111111111001111110010000000000000000;
				player_sprite[840+:120] = 120'b000000000000000011111111111111111111111111111001111110011111100100000000111110010000000011111111000000000000000000000000;
				player_sprite[720+:120] = 120'b000000000000000000000000000000000000000011111001111110011111100111111001111110011111100100000000000000000000000000000000;
				player_sprite[600+:120] = 120'b000000001110000000000000000000001111100111111001111110011111100111111001000000001111100100000000000000000000000000000000;
				player_sprite[480+:120] = 120'b000000000000000000000000010001000100010011111001000000000000000011111001111110010000000000000000000000000000000000000000;
				player_sprite[360+:120] = 120'b000000000000000011100000010001001110000011100000111000001110000011100000111000001110000000000000000000000000000000000000;
				player_sprite[240+:120] = 120'b000000000000000000000000010001000100010011100000111000001110000011100000111000000100010000000000000000000000000000000000;
				player_sprite[120+:120] = 120'b000000000000000000000000000000000100010001000100010001000100010001000100010001000100010000000000000000000000000000000000;
				player_sprite[0+:120] = 120'b000000000000000000000000000000000000000001000100010001000100010001000100010001000000000000000000000000000000000000000000;
			end
			2'd1: begin
				player_sprite[2280+:120] = 120'b111110011111100100000000000000000000000000000000111110011111100111111001000000000000000000000000000000000000000000000000;
				player_sprite[2160+:120] = 120'b111110011111100100000000000000000000000000000000000000001111100111111001000000000000000000000000000000000000000000000000;
				player_sprite[2040+:120] = 120'b000000001111100111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000;
				player_sprite[1920+:120] = 120'b000000001111111111111111010001000000000000000000000000001111100111111111000000000000000000000000000000000000000000000000;
				player_sprite[1800+:120] = 120'b000000000000000011111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000;
				player_sprite[1680+:120] = 120'b000000000000000011111111111111111111111100000000111111111111111100000000000000000000000000000000000000000000000000000000;
				player_sprite[1560+:120] = 120'b000000000000000011111111010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				player_sprite[1440+:120] = 120'b000000000000000000000000111000001110000000000000111111110100010000000000000000000000000000000000000000000000000000000000;
				player_sprite[1320+:120] = 120'b000000000000000011111001111000001110000011111001000000001111111100000000000000000000000000000000000000000000000000000000;
				player_sprite[1200+:120] = 120'b000000000000000011111001111000001110000011100000111110011111100100000000000000000000000000000000000000000000000000000000;
				player_sprite[1080+:120] = 120'b000000000000000011111001010001001111100101000100010001001111100111111001111110011111100111111001000000001111100111100000;
				player_sprite[960+:120] = 120'b000000000000000011111001111110011111100100000000111110011111100100000000111000001111100111111001000000000000000011100000;
				player_sprite[840+:120] = 120'b000000000000000011111001111110011111111100000000111110011111100111111001111110010000000000000000000000001110000011100000;
				player_sprite[720+:120] = 120'b000000000000000000000000000000001111111111111001111110011111100111111001111110010000000000000000000000000000000000000000;
				player_sprite[600+:120] = 120'b000000000000000000000000000000000000000011111001000000001111100111111001111110010000000000000000000000000000000000000000;
				player_sprite[480+:120] = 120'b000000000000000011100000000000000000000000000000000000001111100100000000111110010000000000000000000000000000000000000000;
				player_sprite[360+:120] = 120'b000000000000000000000000111000000000000011100000111000001110000011100000111000000000000000000000000000000000000000000000;
				player_sprite[240+:120] = 120'b000000000000000000000000000000000000000001000100010001000100010001000100010001000100010000000000000000000000000000000000;
				player_sprite[120+:120] = 120'b000000000000000000000000000000000000000001000100010001000100010001000100010001000000000000000000000000000000000000000000;
				player_sprite[0+:120] = 120'b000000000000000000000000000000000000000001000100010001000100010000000000000000000000000000000000000000000000000000000000;
			end
			2'd2: begin
				player_sprite[2280+:120] = 120'b000000001111100111111001111110011111100100000000000000000000000000000000000000001111100111111001111110011111100100000000;
				player_sprite[2160+:120] = 120'b000000001111100111111001111110011111100100000000000000000000000000000000000000001111100111111001111110011111100100000000;
				player_sprite[2040+:120] = 120'b000000000000000011111001111110011111100100000000000000000000000001000100000000001111100111111001000000000000000000000000;
				player_sprite[1920+:120] = 120'b000000000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111000000000000000000000000;
				player_sprite[1800+:120] = 120'b000000000000000011111111111111111111111111111111111111110000000011111111111111111111111111111111000000000100010000000000;
				player_sprite[1680+:120] = 120'b000000000000000000000000111111111111111111111111111111110000000011111111000000001111111111111111000000000000000000000000;
				player_sprite[1560+:120] = 120'b000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
				player_sprite[1440+:120] = 120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				player_sprite[1320+:120] = 120'b000000000000000000000000000000001111100111111001111110011111100100000000111000001110000000000000111110011111100100000000;
				player_sprite[1200+:120] = 120'b000000000000000000000000000000001111100111111001111110010000000000000000111000001110000000000000111110011111100100000000;
				player_sprite[1080+:120] = 120'b000000000000000000000000111111111111100111111001000000001111111100000000111000001110000000000000111110011111100100000000;
				player_sprite[960+:120] = 120'b000000000000000000000000111111111111100111111001000000000000000011111001111110011111111100000000000000000000000000000000;
				player_sprite[840+:120] = 120'b000000000000000000000000000000001111111111111111000000001111100111111001111110010000000000000000111000001110000000000000;
				player_sprite[720+:120] = 120'b000000000000000001000100000000000000000001000100111110011111100111111001111110011111100100000000111000001110000000000000;
				player_sprite[600+:120] = 120'b000000000000000000000000111000000000000011111001000000001111100111111001111110011111100100000000000000001110000000000000;
				player_sprite[480+:120] = 120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				player_sprite[360+:120] = 120'b000000000000000000000000000000000100010000000000010001000100010001000100111000000100010001000100000000000000000000000000;
				player_sprite[240+:120] = 120'b000000000000000000000000000000000000000001000100010001000100010001000100010001000100010001000100010001000000000000000000;
				player_sprite[120+:120] = 120'b000000000000000001000100000000000000000001000100010001000100010001000100010001000100010001000100000000000000000000000000;
				player_sprite[0+:120] = 120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			end
			default: player_sprite = 0;
		endcase
		if (is_1_displayed) begin
			if (~p1Left) begin : sv2v_autoblock_1
				reg signed [31:0] i;
				for (i = 0; i < player_height; i = i + 1)
					begin : sv2v_autoblock_2
						reg signed [31:0] j;
						for (j = 0; j < player_width; j = j + 1)
							player[(((player_height * player_width) * 8) - 1) - (((i * player_width) + j) * 8)-:8] = player_sprite[((i * player_width) + ((player_width - 1) - j)) * 8+:8];
					end
			end
			else begin : sv2v_autoblock_3
				reg signed [31:0] i;
				for (i = (player_height * player_width) - 1; i >= 0; i = i - 1)
					player[(((player_height * player_width) * 8) - 1) - (i * 8)-:8] = player_sprite[i * 8+:8];
			end
		end
		else if (is_2_displayed) begin
			if (~p2Left) begin : sv2v_autoblock_4
				reg signed [31:0] i;
				for (i = (player_height * player_width) - 1; i >= 0; i = i - 1)
					player[(((player_height * player_width) * 8) - 1) - (i * 8)-:8] = player_sprite[i * 8+:8];
			end
			else begin : sv2v_autoblock_5
				reg signed [31:0] i;
				for (i = 0; i < player_height; i = i + 1)
					begin : sv2v_autoblock_6
						reg signed [31:0] j;
						for (j = 0; j < player_width; j = j + 1)
							player[(((player_height * player_width) * 8) - 1) - (((i * player_width) + j) * 8)-:8] = player_sprite[((i * player_width) + ((player_width - 1) - j)) * 8+:8];
					end
			end
		end
		else
			player = 0;
	end
	initial _sv2v_0 = 0;
endmodule
