`default_nettype none
module t03_text_lut (
	alphabet,
	characters
);
	reg _sv2v_0;
	parameter signed [31:0] number_of_chars = 12;
	parameter signed [31:0] character_bits = 72;
	parameter signed [31:0] char_size = 6;
	input wire [(char_size * number_of_chars) - 1:0] alphabet;
	output reg [(number_of_chars * character_bits) - 1:0] characters;
	reg [5:0] bit_select;
	wire [4:0] row_indexing;
	parameter y_length = 8;
	parameter x_length = 9;
	parameter width = x_length * y_length;
	reg [character_bits - 1:0] text;
	always @(*) begin
		if (_sv2v_0)
			;
		begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 1; i <= number_of_chars; i = i + 1)
				begin
					begin : sv2v_autoblock_2
						reg signed [31:0] j;
						for (j = 0; j <= (char_size - 1); j = j + 1)
							bit_select[(char_size - 1) - j] = alphabet[(((char_size * number_of_chars) - 1) - j) - (char_size * (i - 1))];
					end
					case (bit_select)
						6'd0: begin
							text[71:63] = 9'b001110000;
							text[62:54] = 9'b010001000;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b100000100;
							text[35:27] = 9'b111111100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b100000100;
						end
						6'd1: begin
							text[71:63] = 9'b111111000;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b111111000;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b111111000;
						end
						6'd2: begin
							text[71:63] = 9'b001111100;
							text[62:54] = 9'b010000000;
							text[53:45] = 9'b100000000;
							text[44:36] = 9'b100000000;
							text[35:27] = 9'b100000000;
							text[26:18] = 9'b100000000;
							text[17:9] = 9'b010000000;
							text[8:0] = 9'b001111100;
						end
						6'd3: begin
							text[71:63] = 9'b111111000;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b100000100;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b111111000;
						end
						6'd4: begin
							text[71:63] = 9'b111111100;
							text[62:54] = 9'b100000000;
							text[53:45] = 9'b100000000;
							text[44:36] = 9'b111111000;
							text[35:27] = 9'b100000000;
							text[26:18] = 9'b100000000;
							text[17:9] = 9'b100000000;
							text[8:0] = 9'b111111100;
						end
						6'd5: begin
							text[71:63] = 9'b111111100;
							text[62:54] = 9'b100000000;
							text[53:45] = 9'b100000000;
							text[44:36] = 9'b111111000;
							text[35:27] = 9'b100000000;
							text[26:18] = 9'b100000000;
							text[17:9] = 9'b100000000;
							text[8:0] = 9'b100000000;
						end
						6'd6: begin
							text[71:63] = 9'b001111100;
							text[62:54] = 9'b010000000;
							text[53:45] = 9'b100000000;
							text[44:36] = 9'b100011100;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111100;
						end
						6'd7: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b111111100;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b100000100;
						end
						6'd8: begin
							text[71:63] = 9'b011111110;
							text[62:54] = 9'b000110000;
							text[53:45] = 9'b000110000;
							text[44:36] = 9'b000110000;
							text[35:27] = 9'b000110000;
							text[26:18] = 9'b000110000;
							text[17:9] = 9'b000110000;
							text[8:0] = 9'b011111110;
						end
						6'd9: begin
							text[71:63] = 9'b000111110;
							text[62:54] = 9'b000001100;
							text[53:45] = 9'b000001100;
							text[44:36] = 9'b000001100;
							text[35:27] = 9'b000001100;
							text[26:18] = 9'b000001100;
							text[17:9] = 9'b100001100;
							text[8:0] = 9'b011111000;
						end
						6'd10: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b100001000;
							text[53:45] = 9'b100010000;
							text[44:36] = 9'b111100000;
							text[35:27] = 9'b100010000;
							text[26:18] = 9'b100001000;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b100000010;
						end
						6'd11: begin
							text[71:63] = 9'b100000000;
							text[62:54] = 9'b100000000;
							text[53:45] = 9'b100000000;
							text[44:36] = 9'b100000000;
							text[35:27] = 9'b100000000;
							text[26:18] = 9'b100000000;
							text[17:9] = 9'b100000000;
							text[8:0] = 9'b111111100;
						end
						6'd12: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b110001100;
							text[53:45] = 9'b101010100;
							text[44:36] = 9'b100100100;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b100000100;
						end
						6'd13: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b110000100;
							text[53:45] = 9'b101000100;
							text[44:36] = 9'b100100100;
							text[35:27] = 9'b100010100;
							text[26:18] = 9'b100001100;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b100000100;
						end
						6'd14: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b100000010;
							text[44:36] = 9'b100000010;
							text[35:27] = 9'b100000010;
							text[26:18] = 9'b100000010;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111000;
						end
						6'd15: begin
							text[71:63] = 9'b111111000;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b111111000;
							text[35:27] = 9'b100000000;
							text[26:18] = 9'b100000000;
							text[17:9] = 9'b100000000;
							text[8:0] = 9'b100000000;
						end
						6'd16: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b100000010;
							text[44:36] = 9'b100000010;
							text[35:27] = 9'b100000010;
							text[26:18] = 9'b100010010;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111010;
						end
						6'd17: begin
							text[71:63] = 9'b111111000;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b111111000;
							text[35:27] = 9'b100010000;
							text[26:18] = 9'b100001000;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b100000010;
						end
						6'd18: begin
							text[71:63] = 9'b011111100;
							text[62:54] = 9'b100000000;
							text[53:45] = 9'b100000000;
							text[44:36] = 9'b011111000;
							text[35:27] = 9'b000000100;
							text[26:18] = 9'b000000100;
							text[17:9] = 9'b000000100;
							text[8:0] = 9'b111111000;
						end
						6'd19: begin
							text[71:63] = 9'b111111110;
							text[62:54] = 9'b000110000;
							text[53:45] = 9'b000110000;
							text[44:36] = 9'b000110000;
							text[35:27] = 9'b000110000;
							text[26:18] = 9'b000110000;
							text[17:9] = 9'b000110000;
							text[8:0] = 9'b000110000;
						end
						6'd20: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b100000100;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b010001000;
							text[8:0] = 9'b001110000;
						end
						6'd21: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b100000100;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b010001000;
							text[17:9] = 9'b001110000;
							text[8:0] = 9'b000100000;
						end
						6'd22: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b100000100;
							text[53:45] = 9'b100000100;
							text[44:36] = 9'b100100100;
							text[35:27] = 9'b100100100;
							text[26:18] = 9'b101010100;
							text[17:9] = 9'b110001100;
							text[8:0] = 9'b100000100;
						end
						6'd23: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b010001000;
							text[53:45] = 9'b001110000;
							text[44:36] = 9'b000100000;
							text[35:27] = 9'b001110000;
							text[26:18] = 9'b010001000;
							text[17:9] = 9'b100000100;
							text[8:0] = 9'b100000100;
						end
						6'd24: begin
							text[71:63] = 9'b100000100;
							text[62:54] = 9'b010001000;
							text[53:45] = 9'b001110000;
							text[44:36] = 9'b000100000;
							text[35:27] = 9'b000100000;
							text[26:18] = 9'b000100000;
							text[17:9] = 9'b000100000;
							text[8:0] = 9'b000100000;
						end
						6'd25: begin
							text[71:63] = 9'b111111110;
							text[62:54] = 9'b000000100;
							text[53:45] = 9'b000001000;
							text[44:36] = 9'b000010000;
							text[35:27] = 9'b000100000;
							text[26:18] = 9'b001000000;
							text[17:9] = 9'b010000000;
							text[8:0] = 9'b111111110;
						end
						6'd26: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b100001010;
							text[44:36] = 9'b100010010;
							text[35:27] = 9'b100100010;
							text[26:18] = 9'b101000010;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111000;
						end
						6'd27: begin
							text[71:63] = 9'b000110000;
							text[62:54] = 9'b001110000;
							text[53:45] = 9'b000110000;
							text[44:36] = 9'b000110000;
							text[35:27] = 9'b000110000;
							text[26:18] = 9'b000110000;
							text[17:9] = 9'b000110000;
							text[8:0] = 9'b011111110;
						end
						6'd28: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b000000100;
							text[44:36] = 9'b000001000;
							text[35:27] = 9'b000110000;
							text[26:18] = 9'b001000000;
							text[17:9] = 9'b010000000;
							text[8:0] = 9'b011111110;
						end
						6'd29: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b000000100;
							text[44:36] = 9'b000111000;
							text[35:27] = 9'b000000100;
							text[26:18] = 9'b000000100;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111000;
						end
						6'd30: begin
							text[71:63] = 9'b000001000;
							text[62:54] = 9'b000011000;
							text[53:45] = 9'b000101000;
							text[44:36] = 9'b001001000;
							text[35:27] = 9'b010001000;
							text[26:18] = 9'b011111110;
							text[17:9] = 9'b000001000;
							text[8:0] = 9'b000001000;
						end
						6'd31: begin
							text[71:63] = 9'b011111110;
							text[62:54] = 9'b010000000;
							text[53:45] = 9'b010000000;
							text[44:36] = 9'b011111000;
							text[35:27] = 9'b000000100;
							text[26:18] = 9'b000000100;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111000;
						end
						6'd32: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b100000000;
							text[44:36] = 9'b111111000;
							text[35:27] = 9'b100000100;
							text[26:18] = 9'b100000100;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111000;
						end
						6'd33: begin
							text[71:63] = 9'b011111110;
							text[62:54] = 9'b000000100;
							text[53:45] = 9'b000001000;
							text[44:36] = 9'b000010000;
							text[35:27] = 9'b000100000;
							text[26:18] = 9'b001000000;
							text[17:9] = 9'b010000000;
							text[8:0] = 9'b100000000;
						end
						6'd34: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b010000100;
							text[44:36] = 9'b001111000;
							text[35:27] = 9'b010000100;
							text[26:18] = 9'b010000100;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111000;
						end
						6'd35: begin
							text[71:63] = 9'b001111000;
							text[62:54] = 9'b010000100;
							text[53:45] = 9'b010000100;
							text[44:36] = 9'b001111100;
							text[35:27] = 9'b000000100;
							text[26:18] = 9'b000000100;
							text[17:9] = 9'b010000100;
							text[8:0] = 9'b001111000;
						end
						default: text[71:0] = 72'd0;
					endcase
					begin : sv2v_autoblock_3
						integer j;
						for (j = 0; j < y_length; j = j + 1)
							begin : sv2v_autoblock_4
								reg signed [31:0] k;
								for (k = 0; k < x_length; k = k + 1)
									characters[((((number_of_chars * character_bits) - 1) - ((number_of_chars * x_length) * j)) - (x_length * (i - 1))) - k] = text[((character_bits - 1) - (x_length * j)) - k];
							end
					end
				end
		end
	end
	initial _sv2v_0 = 0;
endmodule
